module AFIFO_TEST(
	input rst, clk1,clk2,
	input[7:0] input_data,
	output
	

);

endmodule