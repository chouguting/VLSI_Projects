library verilog;
use verilog.vl_types.all;
entity TESTBED is
end TESTBED;
