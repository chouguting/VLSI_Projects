library verilog;
use verilog.vl_types.all;
entity AFIFO_vlg_vec_tst is
end AFIFO_vlg_vec_tst;
