library verilog;
use verilog.vl_types.all;
entity Lab1Test_vlg_vec_tst is
end Lab1Test_vlg_vec_tst;
