library verilog;
use verilog.vl_types.all;
entity CDC_vlg_vec_tst is
end CDC_vlg_vec_tst;
