library verilog;
use verilog.vl_types.all;
entity Lab1Test_vlg_check_tst is
    port(
        \out\           : in     vl_logic_vector(9 downto 0);
        sampler_rx      : in     vl_logic
    );
end Lab1Test_vlg_check_tst;
